package my_pkg;

  `include "uvm_macros.svh"
   import uvm_pkg ::*;
  `include "transaction.sv"
  `include "sequence.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "agent.sv"
  `include "env.sv"
 // `include "coverage.sv"
endpackage
